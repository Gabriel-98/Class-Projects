LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY TB_alu IS
END TB_alu;
 
ARCHITECTURE behavior OF TB_alu IS 
    COMPONENT alu
    PORT(
         A : IN  std_logic_vector(7 downto 0);
         B : IN  std_logic_vector(7 downto 0);
         C : IN  std_logic_vector(7 downto 0);
         Sc2 : IN  std_logic;
         Sc1 : IN  std_logic;
         Sc0 : IN  std_logic;
         Cout : OUT  std_logic;
         S : OUT  std_logic_vector(7 downto 0)
        );
    END COMPONENT;

   signal A : std_logic_vector(7 downto 0) := (others => '0');
   signal B : std_logic_vector(7 downto 0) := (others => '0');
   signal C : std_logic_vector(7 downto 0) := (others => '0');
   signal Sc2 : std_logic := '0';
   signal Sc1 : std_logic := '0';
   signal Sc0 : std_logic := '0';
   signal Cout : std_logic;
   signal S : std_logic_vector(7 downto 0);
   
BEGIN
   uut: alu PORT MAP (
          A => A,
          B => B,
          C => C,
          Sc2 => Sc2,
          Sc1 => Sc1,
          Sc0 => Sc0,
          Cout => Cout,
          S => S
        );
		  
   stim_proc: process
   begin		
      A <= "00101100";
		B <= "00100110";
		C <= "00110010";
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		A <= "00111100";
		B <= "00011010";
		C <= "00100010";
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		A <= "00001000";
		B <= "00110011";
		C <= "00100101";
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		A <= "00101001";
		B <= "00100110";
		C <= "00100011";
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		A <= "00100110";
		B <= "00101110";
		C <= "00100100";
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		A <= "00110110";
		B <= "00110110";
		C <= "00001100";
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '0';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '0';
		Sc0 <= '1';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '0';
      wait for 20 ns;
		Sc2 <= '1';
		Sc1 <= '1';
		Sc0 <= '1';
      wait for 20 ns;	
   end process;

END;
